`timescale 1ns / 1ps

module processor(clk );


endmodule
